module test (
  input wire a,
  output wire b
);
  
endmodule
