module bnn (
  input wire a,
  input wire b
);
  
endmodule
