module xnor_popcount (
  input wire []
  input wire

  output wire
);
  
endmodule