module shift_reg (
  input wire 
);
  
endmodule